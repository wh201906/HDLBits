module top_module( 
    input [3:0] in,
    output [2:0] out_both,
    output [3:1] out_any,
    output [3:0] out_different );

    always@(*) begin
        casez(in):
            4'b1???:
            
    end

endmodule
