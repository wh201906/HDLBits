module top_module(
    input clk,
    input load,
    input [511:0] data,
    output [511:0] q
);
    wire [511:0] Lq,Rq;
    assign Lq={1'b0,q[511:1]};
    assign Rq={q[510:0],1'b0};
    
    always@(posedge clk) begin
        if(load)
            q<=data;
        else
            q<=~Rq&q | ~Lq&Rq | Lq&~q&Rq;
    end

endmodule
